module pra1 ( 
	a,
	b,
	c,
	d,
	e,
	f,
	g,
	h,
	i,
	j
	) ;

input  a;
input  b;
inout  c;
inout  d;
inout  e;
inout  f;
inout  g;
inout  h;
inout  i;
inout  j;

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SERIES IS
	PORT(
		CLK, CLR: IN STD_LOGIC;
		S: IN STD_LOGIC;
		SHIFTLOAD: IN STD_LOGIC;
		D: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		Q: OUT STD_LOGIC
		);
	ATTRIBUTE PIN_NUMBERS OF SERIES: ENTITY IS "CLK:1, CLR:2, SHIFTLOAD:3, D(3):4, D(2):5, D(1):6, D(0):7";
END ENTITY;

ARCHITECTURE A_SERIES OF SERIES IS
SIGNAL QAUX: STD_LOGIC_VECTOR (3 DOWNTO 0);
BEGIN 
	PROCESS(CLK, CLR) BEGIN
		IF (CLR ='1') THEN
			QAUX <= (OTHERS => '0');
		ELSIF (CLK'EVENT AND CLK = '1') THEN 
			IF (SHIFTLOAD = '1') THEN 
				QAUX <= D;
			ELSE 
				QAUX(2 DOWNTO 0) <= QAUX(3 DOWNTO 1);
				QAUX(3) <= S;
			END IF;
		END IF;
	END PROCESS;
	Q <= QAUX(0);
END A_SERIES;

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SERIES IS
	PORT(
		CLK, CLR: IN STD_LOGIC;
		D: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		Q: OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
		);

END ENTITY;

ARCHITECTURE A_SERIES OF SERIES IS
SIGNAL Q1, Q2: STD_LOGIC;
BEGIN 
	PROCESS(CLK, CLR) BEGIN
		IF (CLR ='1') THEN
			Q <= (OTHERS => '0');
		ELSIF (CLK'EVENT AND CLK = '1') THEN 
			Q<= D;
		END IF;
	END PROCESS;
END A_SERIES;
module series ( 
	clk,
	clr,
	d,
	q
	) ;

input  clk;
input  clr;
input [3:0] d;
inout [3:0] q;

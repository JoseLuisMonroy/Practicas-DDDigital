module series ( 
	d,
	clk,
	clr,
	q
	) ;

input  d;
input  clk;
input  clr;
inout  q;

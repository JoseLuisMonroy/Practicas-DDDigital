LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY DETECTOR IS 
	PORT( CLK :IN STD_LOGIC;
	CLR: IN STD_LOGIC;
	ENTRADA: IN STD_LOGIC;
	SALIDA: OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
END DETECTOR;

ARCHITECTURE COMPORTAMENTAL OF DETECTOR IS 
TYPE ESTADOS IS(A, B, C, D, E, F, G);		  
attribute ENUM_ENCODING: STRING;
ATTRIBUTE enum_encoding OF ESTADOS: TYPE IS
"0000" & --A--	  
"0001" & --B--
"0011" & --C--
"0010" & --D--
"0110" & --E--
"0111" & --F--
"1111" ; --G--
SIGNAL EDO, NEXT_EDO: ESTADOS; 
BEGIN

PROCESS (CLR, CLK)
BEGIN 
	IF(CLR = '1') THEN
		EDO <= A;
	ELSIF(CLK'EVENT AND CLK = '1') THEN
		EDO <= NEXT_EDO;
	END IF;
END PROCESS;

PROCESS (ENTRADA, EDO)
BEGIN 
	CASE EDO IS WHEN 
		A => IF ENTRADA = '0' THEN
			NEXT_EDO <= C;
		ELSIF ENTRADA = '1' THEN
			NEXT_EDO <= B;
		END IF;
		WHEN
		B => IF ENTRADA = '0' THEN 
			NEXT_EDO <= C;
		ELSIF ENTRADA = '1' THEN
			NEXT_EDO  <= F;
		END IF;	
		WHEN
		C => IF ENTRADA = '0' THEN 
			NEXT_EDO <= D;
		ELSIF ENTRADA ='1' THEN
			NEXT_EDO <= B;
		END IF;
		WHEN
		D => IF ENTRADA = '0' THEN 
			NEXT_EDO <= E;
		ELSIF ENTRADA ='1' THEN
			NEXT_EDO <= B;
		END IF;			 
		WHEN
		E => IF ENTRADA = '0' THEN 
			NEXT_EDO <= E;
		ELSIF ENTRADA ='1' THEN
			NEXT_EDO <= B;
		END IF;			  
		WHEN
		F => IF ENTRADA = '0' THEN 
			NEXT_EDO <= C;
		ELSIF ENTRADA ='1' THEN
			NEXT_EDO <= G;
		END IF;			  
		WHEN
		G => IF ENTRADA = '0' THEN 
			NEXT_EDO <= C;
		ELSIF ENTRADA ='1' THEN
			NEXT_EDO <= G;
		END IF;		   
		WHEN OTHERS => NULL;
	END CASE;
END PROCESS;
--A B C D E F G--
SALIDA <= "0110000" WHEN (EDO = C AND ENTRADA = '0') ELSE--A--
	"0110000" WHEN (EDO = B AND ENTRADA = '1' ) ELSE 
	"0110000" WHEN (EDO = C AND ENTRADA = '0') ELSE --B--
	"0110000" WHEN (EDO = F AND ENTRADA = '1' ) ELSE
	"0110000" WHEN (EDO = D AND ENTRADA = '0') ELSE --C--
	"0110000" WHEN (EDO = B AND ENTRADA = '1' ) ELSE
	"0001001" WHEN (EDO = E AND ENTRADA = '0') ELSE	--D--
	"0110000" WHEN (EDO = B AND ENTRADA = '1' ) ELSE 
	"0001001" WHEN (EDO = E AND ENTRADA = '0') ELSE	 --E-
	"0110000" WHEN (EDO = B AND ENTRADA = '1' ) ELSE
	"0110000" WHEN (EDO = C AND ENTRADA = '0') ELSE	--F--
	"0001001" WHEN (EDO = G AND ENTRADA = '1' ) ELSE
	"0110000" WHEN (EDO = B AND ENTRADA = '0') ELSE	--G
	"0001001" WHEN (EDO = G AND ENTRADA = '1' ) ELSE   
	"0110000";
END COMPORTAMENTAL;
		
	

		
		


module restador ( 
	ci,
	a,
	b,
	cf,
	s
	) ;

input  ci;
input [3:0] a;
input [3:0] b;
inout  cf;
input [3:0] s;

ARCHITECTURE ARQ_FLIPFLOP OF FLIPFLOP IS
SIGNAL CLK_AUX: STD_LOGIC;
SIGNAL CONTADOR: INTEGER RANGE 0 TO 27000000 := 0;
BEGIN 
	
	DIVISOR_FRECUENCIA: PROCESS (CLR, CLK) BEGIN
		IF (CLR= '1') THEN
			CLK_AUX <= '0';
			CONTADOR <= 0;
		ELSIF RISING_EDGE(CLK) THEN
			IF(CONTADOR = 27000000) THEN
				CLK_AUX <= NOT (CLK_AUX);
				CONTADOR <= 0;
			ELSE
				CONTADOR <= CONTADOR + 1;
			END IF;
		END IF;
	END PROCESS;
	SALIDA <= CLK_AUX; 
END ARQ_FLIFLOP;

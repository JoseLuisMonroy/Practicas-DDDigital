LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY PR1 IS

PORT(
	A: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	F: OUT STD_LOGIC
	);

ATTRIBUTE PIN_NUMBERS OF PR1:ENTITY IS "A(0):1 A(1):2 A(2):3 A(3):4 F:17";

END ENTITY;

ARCHITECTURE A_PR1 OF PR1 IS

BEGIN
	F <= ((A(0) AND A(1))AND (NOT A(2)))OR ((A(1) AND A(2))AND A(3));

END ARCHITECTURE;

module series ( 
	d,
	clk,
	clr,
	q,
	q1,
	q2
	) ;

input  d;
input  clk;
input  clr;
inout  q;
inout  q1;
inout  q2;

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SERIES IS
	PORT(
		CLK, CLR: IN STD_LOGIC;
		SI, SD: IN STD_LOGIC;
		SEL: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		D: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		Q: INOUT STD_LOGIC_VECTOR (3 DOWNTO 0)
		);
	--ATTRIBUTE PIN_NUMBERS OF SERIES: ENTITY IS "CLK:1, CLR:2,D(3):3, D(2):4, D(1):5, D(0):6, SEL(1):7, SEL(0):8, SI:9, SD:10, Q(3):21, Q(2):22, Q(1):20, Q(0):19";
END ENTITY;

ARCHITECTURE A_SERIES OF SERIES IS
BEGIN 
	PROCESS(CLK, CLR) BEGIN
		IF (CLR ='1') THEN
			Q <= (OTHERS => '0');
		ELSIF (CLK'EVENT AND CLK = '1') THEN 
			IF (SEL = "11") THEN 
				Q <= D;
			ELSIF (SEL = "01") THEN 
				Q(2 DOWNTO 0) <= Q(3 DOWNTO 1);
				Q(3) <= SI;
			ELSIF (SEL = "10") THEN
				Q(3 DOWNTO 1) <= Q(2 DOWNTO 0);
				Q(0) <= SD;
			END IF;
		END IF;
	END PROCESS;
END A_SERIES;

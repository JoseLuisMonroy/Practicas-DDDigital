LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SERIES IS
	PORT(
		CLK, CLR: IN STD_LOGIC;
		SEL: IN STD_LOGIC;
		Q: INOUT STD_LOGIC_VECTOR (7 DOWNTO 0)
		);
	--ATTRIBUTE PIN_NUMBERS OF SERIES: ENTITY IS "CLK:1, CLR:2,D(3):3, D(2):4, D(1):5, D(0):6, SEL(1):7, SEL(0):8, ";
END ENTITY;

ARCHITECTURE A_SERIES OF SERIES IS
BEGIN 
	PROCESS(CLK, CLR) BEGIN
		IF (CLR ='1') THEN
			Q <= '0';
		ELSIF (CLK'EVENT AND CLK = '1') THEN 
			IF (SEL = '0') THEN 
				
			ELSE
				
			END IF;
		END IF;
	END PROCESS;
END A_SERIES;
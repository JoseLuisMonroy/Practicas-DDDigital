module pr1 ( 
	a,
	f
	) ;

input [3:0] a;
inout  f;

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY DISPMULT IS 
	PORT( 
	--CLK :IN STD_LOGIC;
	CLR: IN STD_LOGIC;						
	AUX_CLK1: IN STD_LOGIC;
	AUX_CLK: IN STD_LOGIC;
	AN: INOUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	SALIDA: OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
END DISPMULT; 

ARCHITECTURE COMPORTAMENTAL OF DISPMULT IS 	 

CONSTANT H: STD_LOGIC_VECTOR(6 DOWNTO 0):= "1001000";
CONSTANT O: STD_LOGIC_VECTOR(6 DOWNTO 0):= "0000001";
CONSTANT L: STD_LOGIC_VECTOR(6 DOWNTO 0):= "1110001"; 
CONSTANT A: STD_LOGIC_VECTOR(6 DOWNTO 0):= "0001000";	   
CONSTANT G: STD_LOGIC_VECTOR(6 DOWNTO 0):= "1111110"; 
CONSTANT I: STD_LOGIC_VECTOR(6 DOWNTO 0):= "1001111";
CONSTANT P: STD_LOGIC_VECTOR(6 DOWNTO 0):= "0011000"; 
CONSTANT N: STD_LOGIC_VECTOR(6 DOWNTO 0):= "1101010";


TYPE ESTADOS IS(Q0, Q1, Q2, Q3, Q4, Q5, Q6, Q7, Q8, Q9, Q10, Q11, Q12, Q13, Q14, Q15, Q16, Q17, Q18, Q19, Q20, Q21, Q22, Q23, Q24, Q25, Q26, Q27, Q28, Q29, Q30, Q31, Q32);
SIGNAL EDO, NEXT_EDO: ESTADOS;
SIGNAL CONTADORBIN: STD_LOGIC_VECTOR(3 DOWNTO 0):="0000" ;

--SIGNAL AUX_CLK: STD_LOGIC;
--SIGNAL CONTADOR: INTEGER RANGE 0 TO 50000000 := 0; 
--SIGNAL CONTADOR1: INTEGER RANGE 0 TO 50000000 := 0; 
BEGIN 
--	DIVISOR_FRECUENCIA: PROCESS (CLR, CLK) BEGIN
--		IF (CLR= '1') THEN
--			AUX_CLK <= '0';
--			CONTADOR <= 0;
--		ELSIF RISING_EDGE(CLK) THEN
--			IF(CONTADOR = 50000000) THEN
--				AUX_CLK <= NOT (AUX_CLK);
--				CONTADOR <= 0;
--			ELSE
--				CONTADOR <= CONTADOR + 1;
--			END IF;
--		END IF;
--	END PROCESS;	 

--	DIVISOR_FRECUENCIA1: PROCESS (CLR, CLK) BEGIN
--		IF (CLR= '1') THEN
--			AUX_CLK1 <= '0';
--			CONTADOR <= 0;
--		ELSIF RISING_EDGE(CLK) THEN
--			IF(CONTADOR = 50000000) THEN
--				AUX_CLK1 <= NOT (AUX_CLK1);
--				CONTADOR <= 0;
--			ELSE
--				CONTADOR1 <= CONTADOR1 + 1;
--			END IF;
--		END IF;
--	END PROCESS;  

CONTADOR_BINARIO: PROCESS (CLR, AUX_CLK1)
BEGIN
	IF (CLR ='1') THEN
		CONTADORBIN <= "0000"; 
	ELSIF (AUX_CLK1'EVENT AND AUX_CLK1 = '1') THEN
		CONTADORBIN <= CONTADORBIN + 1;
	END IF;
END PROCESS;
	

LOGICA_ENTRADA: PROCESS(CLR, AUX_CLK)
BEGIN
	IF (CLR ='1') THEN
		AN <= "0001"; 
		EDO <= A;
	ELSIF (AUX_CLK'EVENT AND AUX_CLK = '1') THEN 
		EDO <= NEXT_EDO;
		AN(3 DOWNTO 1) <= AN(2 DOWNTO 0);
		AN(0) <= AN(3);
	END IF;
END PROCESS;

MAQUINA: PROCESS (EDO, CONTADORBIN)
BEGIN 
	CASE EDO IS WHEN 
		Q0 => IF CONTADORBIN = "0001" THEN
			NEXT_EDO <= Q1;
		END IF;
		WHEN
		Q1 => IF CONTADORBIN = "0010" THEN
			NEXT_EDO <= Q2;
		END IF;
		WHEN 
		Q2 => IF CONTADORBIN = "0010" THEN
			NEXT_EDO <= Q3;
		ELSIF CONTADORBIN = "0011" THEN
			NEXT_EDO <= Q4; 
		END IF;
		WHEN 
		Q3 => IF CONTADORBIN = "0010" THEN
			NEXT_EDO <= Q2;
		ELSIF CONTADORBIN = "0011" THEN
			NEXT_EDO <= Q4;
		END IF;
		WHEN 
		Q4 => IF CONTADORBIN = "0011" THEN
			NEXT_EDO <= Q5;
		ELSIF CONTADORBIN = "0100" THEN
			NEXT_EDO <= Q7;
		END IF;
		WHEN 
		Q5 => IF CONTADORBIN = "0011" THEN
			NEXT_EDO <= Q6;
		ELSIF CONTADORBIN = "0100" THEN
			NEXT_EDO <= Q7;
		END IF;
		Q6 => IF CONTADORBIN = "0011" THEN
			NEXT_EDO <= Q4;
		ELSIF CONTADORBIN = "0100" THEN
			NEXT_EDO <= Q7;
		END IF;	
		WHEN
		Q7 => IF CONTADORBIN = "0100" THEN
			NEXT_EDO <= Q8;
		ELSIF CONTADORBIN = "0101" THEN
			NEXT_EDO <= Q11;
		END IF;
		WHEN
		Q8 => IF CONTADORBIN = "0100" THEN
			NEXT_EDO <= Q9;
		ELSIF CONTADORBIN = "0101" THEN
			NEXT_EDO <= Q11;
		END IF;				
		WHEN
		Q9 => IF CONTADORBIN = "0100" THEN
			NEXT_EDO <= Q10;
		ELSIF CONTADORBIN = "0101" THEN
			NEXT_EDO <= Q11;
		END IF;			   
		WHEN
		Q10 => IF CONTADORBIN = "0100" THEN
			NEXT_EDO <= Q7;
		ELSIF CONTADORBIN = "0101" THEN
			NEXT_EDO <= Q11;
		END IF;	
		WHEN
		Q11 => IF CONTADORBIN = "0101" THEN
			NEXT_EDO <= Q12;
		ELSIF CONTADORBIN = "0110" THEN
			NEXT_EDO <= Q15;
		END IF;	
		WHEN
		Q12 => IF CONTADORBIN = "0101" THEN
			NEXT_EDO <= Q13;
		ELSIF CONTADORBIN = "0110" THEN
			NEXT_EDO <= Q15;
		END IF;
		WHEN
		Q13 => IF CONTADORBIN = "0101" THEN
			NEXT_EDO <= Q14;
		ELSIF CONTADORBIN = "0110" THEN
			NEXT_EDO <= Q15;
		END IF;	
		WHEN
		Q14 => IF CONTADORBIN = "0101" THEN
			NEXT_EDO <= Q11;
		ELSIF CONTADORBIN = "0110" THEN
			NEXT_EDO <= Q15;
		END IF;	   
		WHEN
		Q15 => IF CONTADORBIN = "0110" THEN
			NEXT_EDO <= Q16;
		ELSIF CONTADORBIN = "0111" THEN
			NEXT_EDO <= Q19;
		END IF;	
		WHEN
		Q16 => IF CONTADORBIN = "0110" THEN
			NEXT_EDO <= Q17;
		ELSIF CONTADORBIN = "0111" THEN
			NEXT_EDO <= Q19;
		END IF;	  
		WHEN
		Q17 => IF CONTADORBIN = "0110" THEN
			NEXT_EDO <= Q18;
		ELSIF CONTADORBIN = "0111" THEN
			NEXT_EDO <= Q19;
		END IF;
		WHEN
		Q18 => IF CONTADORBIN = "0110" THEN
			NEXT_EDO <= Q15;
		ELSIF CONTADORBIN = "0111" THEN
			NEXT_EDO <= Q19;
		END IF;	  
		WHEN
		Q19 => IF CONTADORBIN = "0111" THEN
			NEXT_EDO <= Q20;
		ELSIF CONTADORBIN = "1000" THEN
			NEXT_EDO <= Q23;
		END IF;	
		WHEN
		Q20 => IF CONTADORBIN = "0111" THEN
			NEXT_EDO <= Q21;
		ELSIF CONTADORBIN = "1000" THEN
			NEXT_EDO <= Q23;
		END IF;	   
		WHEN
		Q21 => IF CONTADORBIN = "0111" THEN
			NEXT_EDO <= Q22;
		ELSIF CONTADORBIN = "1000" THEN
			NEXT_EDO <= Q23;
		END IF;	  
		WHEN
		Q22 => IF CONTADORBIN = "0111" THEN
			NEXT_EDO <= Q19;
		ELSIF CONTADORBIN = "1000" THEN
			NEXT_EDO <= Q23;
		END IF;	  
		WHEN
		Q23 => IF CONTADORBIN = "1000" THEN
			NEXT_EDO <= Q24;
		ELSIF CONTADORBIN = "1001" THEN
			NEXT_EDO <= Q27;
		END IF;
		Q24 => IF CONTADORBIN = "1000" THEN
			NEXT_EDO <= Q25;
		ELSIF CONTADORBIN = "1001" THEN
			NEXT_EDO <= Q27;
		END IF;
		Q25 => IF CONTADORBIN = "1000" THEN
			NEXT_EDO <= Q26;
		ELSIF CONTADORBIN = "1001" THEN
			NEXT_EDO <= Q27;
		END IF;	
		Q26 => IF CONTADORBIN = "1000" THEN
			NEXT_EDO <= Q23;
		ELSIF CONTADORBIN = "1001" THEN
			NEXT_EDO <= Q27;
		END IF;
		WHEN
		Q27 => IF CONTADORBIN = "1001" THEN
			NEXT_EDO <= Q28;
		ELSIF CONTADORBIN = "1010" THEN
			NEXT_EDO <= Q30;
		END IF;
		WHEN
		Q28 => IF CONTADORBIN = "1001" THEN
			NEXT_EDO <= Q29;
		ELSIF CONTADORBIN = "1010" THEN
			NEXT_EDO <= Q30;
		END IF;	  
		WHEN
		Q29 => IF CONTADORBIN = "1001" THEN
			NEXT_EDO <= Q27;
		ELSIF CONTADORBIN = "1010" THEN
			NEXT_EDO <= Q30;
		END IF;	
		WHEN
		Q30 => IF CONTADORBIN = "1010" THEN
			NEXT_EDO <= Q31;
		ELSIF CONTADORBIN = "1011" THEN
			NEXT_EDO <= Q32;
		END IF;			  
		WHEN
		Q31 => IF CONTADORBIN = "1010" THEN
			NEXT_EDO <= Q30;
		ELSIF CONTADORBIN = "1011" THEN
			NEXT_EDO <= Q32;
		END IF;
		WHEN
		Q32 => IF CONTADORBIN = "1100" THEN
			NEXT_EDO <= Q0;
		WHEN OTHERS => NULL;
	END CASE;
END PROCESS;

SALIDA <= 
	H WHEN (EDO = Q1 OR EDO = Q2 OR EDO = Q4 OR EDO = Q7 ) ELSE
	O WHEN (EDO = Q3 OR EDO = Q5 OR EDO = Q8 OR EDO = Q14) ELSE
	L WHEN (EDO = Q6 OR EDO = Q9 OR EDO = Q13 OR EDO = Q18) ELSE	 
	A WHEN (EDO = Q10 OR EDO = Q12 OR EDO = Q17 OR EDO = Q22) ELSE
	G WHEN (EDO = Q11 OR EDO = Q16 OR EDO = Q21 OR EDO = Q26) ELSE
	I WHEN (EDO = Q15 OR EDO = Q20 OR EDO = Q25 OR EDO = Q29) ELSE
	P WHEN (EDO = Q19 OR EDO = Q24 OR EDO = Q28 OR EDO = Q31) ELSE
	N WHEN (EDO = Q23 OR EDO = Q27 OR EDO = Q30 OR EDO = Q32) ELSE
	"1111111";
END COMPORTAMENTAL;

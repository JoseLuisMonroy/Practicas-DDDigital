LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY SUMADOR IS
	PORT ( CI: IN STD_LOGIC;
			A,B: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			CF: OUT STD_LOGIC;
			S: IN STD_LOGIC_VECTOR(3 DOWNTO 0)
			);
	END ENTITY;
ARCHITECTURE A_SUMADOR OF SUMADOR IS
	SIGNAL C: STD_LOGIC_VECTOR(0 TO 4);
	BEGIN 
		C(0)<=CI;
		CICLO_1: FOR I IN 0 TO 3 GENERATE
			B(I)<= B(I)XNOR CI;
			S(I)<= A(I) XOR B(I)XOR C(I);
			C(I+1)<=(A(I) AND B(I))OR(A(I)AND C(I))OR (B(I)AND C(I));
		END GENERATE;
		CF <=C(4);
    END A_SUMADOR;
   	
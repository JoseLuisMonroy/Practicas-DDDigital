LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY DETECTOR IS 
	PORT( 
	CLK :IN STD_LOGIC;
	CLR: IN STD_LOGIC;						
	AUX_CLK: INOUT STD_LOGIC;
	AN: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	SALIDA: OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
END DETECTOR; 

